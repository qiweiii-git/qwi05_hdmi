//*****************************************************************************
// Define.vh.
//
// Change History:
//  VER.   Author         DATE              Change Description
//  1.0    Qiwei Wu       Apr. 11, 2020     Initial Release
//*****************************************************************************

`include "Qwi05RegDef.vh"
`include "Qwi05FmtDef.vh"
`include "Qwi05RgbDef.vh"